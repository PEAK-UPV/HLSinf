//
// This file is the header for all files with module defines
//

